module pop_count_parallel(
	input clk, 
	input rst, 
	input [9:0]input_number,
	input start,
	output reg [7:0]count,
	output reg done
);



endmodule
