module pop_count_sequential(
	input clk, 
	input rst, 
	input [9:0]input_number,
	input start,
	output reg [7:0]count,
	output reg done
);



endmodule
